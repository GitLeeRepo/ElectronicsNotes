eNrtXetT4sgW/1dSfLm6g9qPJASr/MAI66VG0BsQd2q9ZSHGMbVI3AR2Zu6U//vtR5JOIAmvBKO2
HyJ0+kWfX5/T5/Tp078qPftpNh5ObWdy6TrPlju1La9y/KvSu261Lm8b3cb51167R1Pa3V6/0T1t
3fa/XrYqx5VKtXJ50e72e/xz+PqyYTY6rX7L5Om8ola36RdxvltuYzIc//Rs0tDUnVlBHlLe7EcL
sYTbq267P9dElzQQr73x+bxFWngYjj0r0mZY+OWlWrm2Xf7bYK0OsA7oPxUAmvLgOk9fK8cksVqZ
On9Ujum7KksOv0wdkoPkJzVpNYAAoE8cLU7S/OLkVViafWaFSW5SWNVoscXCOKkwyRwrTN5hDHSV
PqMdDwuTVwkt46AwqgFeRbTlWna3eWHDABoE9KlFC5M0vzB5FRZmn1lhkpsUrqlAw8AA9BktHHbb
AKJwTQ0Ls5ZhDVI6LZJLBSnkgnFyQdUA2AA0nfyLDpshKoCRCtSw+yQHJ5mm04Ejz2j39WySkfdB
93nrZLCi3U9pXXSf5Ket14GGAHnqsV9P0vziauTHqyFU9dhvJ/9UmPLbVSPxt6usdUIZDCjp5hAH
kkhngDhoSG844shzKeJE18l7jjhoUMQhFC0MjWzEkdykcB3R0SZPHSfDtY5E4ToKBw37hUkr5IlB
csvJhTEfcQMz7kL+qUYKdzFwZMQNHI44QxskGXEN0H9zJAuHDbK6ggr8ikOScaiQoY0DRgfZo84B
UyNDplN66zGs63riVBUDp/uFMU4AC84u7HMYQLkqfaJkrpqMNE5vDtMFkgmYRkkWgWk4SQgyIGFW
8Skq4ELfJU0SPkV91uJzqhU4zDyL4sSiT305yQRr5qPOh2xhoiCUOFHmBo7yNsJdtHneJriLlsHb
KFvRgD9+Ud6mLeMuWsBdfMGgLRcMoutcqhDowjrgPCY6TevZjJFzF396LTJGFSZ3fX6W8U4vCkQt
e9R51yEhuz9wqrbSwIUVqIFE9ScLWD5ZhERFICqSFlhURCTFWFQErob/2wmnXOCuOs6ebXqwDCG4
JQuVNA6TvIbhWKeDVgd8DZVMcy1z9aThBDmOs2eZj3XSe8okFuR4hEnE5riO41jnrZOfkbYI0vXE
1rFYcpIcafROLuzTm6CHShQOumSJooIMtHF6LwqFJdOUkoyUPnWenp2JNZl6A9v6TpbjvdGj9USU
jhFd1E+86XAy4ivzwf0Ikve/bioPY/v5pnJ8U/lE/m4q1ZvKKKilO3yy2Kv70cHAGU+H36yDnjNz
RxbL9xzqMSzTn79ubm4qg8b5VYt+OKYPnT6q9NE7bzdbptn6z1XbbDXDDEyPCDN1G/32gGsdYY4r
UcVl67TdOGeqRjxPmKXZ6p2a7ct++6IbvvyH91yxJwr9EV6kteXNxH+OyPPvi+vbS/PismX2v4av
qY4lslx9Pm2bp1fplfy73Wy2uilDEetFs/V74+q8n/B7rzqXVCNb2oXk4eq0u3OdA0mF25xek9l4
zF4tEmBQfRpUZ4OwcMLYVa0DgOlDYKLT+CO1ear7hslmq3Eer3t+RFjBl/8yXFLt9bb3tfP54pwB
8/fx0HtsnvoIZlm8n093zvjS8WyqkJNcZCL8JP80wpZvKj9u2Mx+qcYRSesi84ZV4DrToV/0pgIh
S4uCj88aJcCeJ2ZNQqNa7VALmlXRoUYbPm9/Nhvm19sz8+LqklUXn5u305/PfHIOiY7vfGNvbX+K
hxOXTnP2hg1n9Aect09b3R63MbAXgA+MNbZGU+v+Mj63r9jLVrPdZ2ijSQxprMjsrml5I9d+Dgfk
SjlRdIXAYcIHiwzV5BtnEoREL5QZdayp5c6zoIODVBbUeHqiJRIZTwbZo8XSiE4ZOh993UgkepuM
xp21SHcAEukebTOhNbUetIZzpLQ/oHFi88QseieTNIFgzU5HW11gNO1v9nQ4PujMxlObjcYBgv5w
zVGPSY2riT0N5zIEiuAkzIwlXgn2xGZUnw5NyISap4wLZDCBTifsRhoasBqgAeJkOJBaVsaCPxCK
GAgl7EFC20AL29ZAfuCgxIsjI/gNC7CA68Gib/2YQrQ6MGj+g8ZkEg5d2joixv/7rT/66fw/lEtx
WeLze+ViNlXogomk3UyCxKb9j33PgHUzaf09452hXw4W/3hBe3KiD9hHE5/ALxePvEJTPUHhl0Hz
xFSP9kz8yVT3gxR0hP2mZ9OTQfM3UpP4jgfbr5CGYjiz1kF81EkuhRIheRWUUNVqC5GlS43kFdPc
mme7JdPCYij+OnOxs3xpudZ6aKUlzioLzZR3WSsdSt25GZYq+QSvAyiR1yVUtpIIvL8nnIIDLUUM
4qDpei1HTsf5UZzXhb1Yb82z3pInjUGS9RaQipZUtKSiFZv+SHsFRQuhIhUtUEpFy1zDzGNanu1N
HXdVpgO3ZzrmtkyH95nSIpndmJLdbMFuyMLWq35hzw59ZvOdT5TvfCqG7zCsvVQTUIj0Q0PbHol9
6+l5WzB6oY+HMiXVWWQ+zlwmEO+tb65lKafWeGTPUiRjeg/WQuuWa+o40t4UWpetmvPGZCokQQ5w
HMFt0fhgu95UcVyi58bgOHKshwd7ZBPWnwLEtLYlDj8gDtHWXNEaOZP7zYCIJBDfAxDzktETZsbb
Co1RAA6nyvdHe/SoPA/dIbPOesp3i7ywfkzdIV2ep+AytR8SmOUFZobSGtN8UnVWEOisNZCos5or
28fOrInl2iMl1u5ii9TZwt8r0tQ81VVzbqPI3EBVNddTVU2iqkLlC9ciFtXVJOl1iDSwqnU3iV1k
8oHO8AdZrT8pd641/Et5pttMynDkOp6nuD5VDpNn/yUpGodb7PXTdfW6+uV6BXUmbQYwAw5TpzIY
SDi7YlMh3C7L1ERfors3uNS7N/5GjTLzqEGZU4ayaaJT9cgUsrxtACJ3TtYQyHL/ZNFzA4r9E2O3
+ycaEE3jvDdQcIk2UJqdDvwQjgcwNInXwY79DiAMzOJGLV+3A1ig24FWSsHVd+i4x8zSNxOzf6KY
8JOJ2LfrR6pjmH3F9pSE7Ms53yvIsnTu/WEE2EriPEsbzV6glMAdYJnnU4HSLGw5d2GmlUuY4Q8h
zNRQc1VrOxZmqhYIM1XNV5jhYoTZAA1Xx8T58M4ar+sFSw/kioKpC5CQZoaaSLOVCdZ17i1FNJjQ
VA0fijUHxLluxaNhnE6iI9tOec6wE+c8F4fJ5L0rBXnpQbMdkVcDRZL3rlTkPZvcr+H/euY6s8n9
ugSOlFpOXagmC+8zv4aV7JOiwSTqhl7KqmbkSVs6lnHiBp3e1n2drQSMUioMpzPX5Ttgce/j1d2O
iXbBXI6DLzh80z4hFRyZff+L7rsit09Qp8GcDehncAgAakg/ZOmHXAI/ZPhqfsgQ5O6IbJRI9TC1
PB0BN/HeqhbsQZije2De/CVPD8LsPdxdcpdU78ACuE3cu9B3MthgF7i6GwfCXXoHlkwYxuBYHrAW
LgrzhGTODoS78Q6UOJQ4zHYg3JF3oATiuwNiEQ6Eu/cOlMAsu9K6kiOgKtTVGlzVEzDl7NqKnoCq
UFN1PV9XQK2UroCbObytpXy+E//CTGVxqXdh1BUQLZ5UPjgoVyAHZrKk0RwUgp5/ecr58Htm2Aaz
H7GTtk9waPZk0Rfae2Z/X3xFe4cA4P3E6AzSHUO6Y+zYKorC/ViI8G6tosgQBlkjZ6soAmWyiqol
tIqijblObsbQ3PnL27GAbshXUo2hKzHDsltF1wXiTo2hZROGO9SrthWCRYKzQGvU2nDciTFU4lDi
EJTBGCqB+DGAuKWM3r0xVAKzvMDc1iqqCfdhsBujqIjWXMv5eLT6KjZRJG2ipbKJNjsd9WPEPBa7
Cwbc8XENVA+9iWtGvuc11AIPH4JS+hL37KfnMdGdbXc0s4nEtqePCvTZaIQlSBdf6eK7Y2M2FocL
6/XdGrOxOF1YV/N28S2TMZt1SC0lY4rv1rVPBkcm32Y7afMPJklqy902udv2WgyqJjbbtB0fQRAt
g7zZk1oi9nQ2uYclOCmn15aEns7toJyuiWjTeZ+Tg8Wck+M3xqBS3MsTia6j1Yu/mEet18Pm1Nxv
5kGF3cxDSA9KMK3EvTlFTyuMiptWoJhpRZXwjxH3wXi1IEaqWlQQI1SgHaH+ps4kLx5K1qKHkvsn
phZ8gumHkGHwae4Qsi4PIUsLxaspACJkDQI71gAE1yQaQN4qQL1ctyEheRuSvA1J3oaUdrojJXhL
EdchqUBchwRVLe/7kFAp70NiLFF/EyGPY/dSsvMIJjraY2Ek9/fIkmpfrpbkaum1VktQxJvCtd2u
lqCwC2GU92pJL9PhBFTqkC3ZqwAZq6WMgdXfZciW9YEoY7UkYf3D3QJQjFP4BnCUsVokDkuBQxmr
RQKxLDJaxmqRwMzt7jZ914cTxA3neR9OQDJgizycwCwTRqntmDReCw3V4tsvY8ZNlhYYOJW91t/K
d8f9y2PJ1j8W0boendm3R/KPMHGWanvKxFGCaliSX9d+ZgSYtM3qQfPE1I78/WryBQoz66AZmFf9
BF3GgZGeqa93yxya91/f3b08wtRq1HM2tRrlupcHfIxL5vRXu5cHoqLu5QHF+Wfh9yFhV5aQMOrO
hebEZbj7GMrMIxSVmr+RmhKDp8mrWeXVrLs+b4bm70fd3XmzUGjW846dhst22qz2tq/USWV31JU1
vK9zLojknDcrWogtyb1ZcUMqDSX0xXjLcTg243/w1fhfcCt2jv4ZtZJxQATfY8zc6A1iKDNmLqYx
c9G+XPbJZV8pbhKDrxYzVwcFxsyFZXLiR6NSXGiKxZHtmlbwjaZYi9xoCmso5ytNR6W60pQhDpVy
Zd91ppYyfRxO6c6AYvnmDb5vMPMstkelPDiuYvaV4eSepRPx5bE0Xy1Q9trSdVq6Tr+e67QIro53
fNAMCpaJ8z5ohlCZXKdxnq7TBV5aueHpsg19peW5su28pJd6Oed9wAxG3LKKv7VyQzAW5Sy9Flpz
9a96U2hdJrbyxmQqJHO+tXJDNObvLC1x+AFxiLbmivk7S0sgvi0gFnFr5YZoLNZZWgKzvMDcOq57
GJygtrLrdFpYrxXjuod7V3rOrtO4lK7T79LLeYln91I/5+rmTuVpmuhLLMghKEWQQxF6XTeKj3GI
YRDjUMe5hzgEhYU4pKYk8CZidsw8aoFz/YDrHtWBe4TlWZ7cFJWboiUwOAPj1QzOvhtefgbn8oRe
f6lW/uc4T/RHgmolcLr1Ksd//qo825O+c+ba94R/AcLL4kQiiagOfiBAaP3yfxUgpNY=