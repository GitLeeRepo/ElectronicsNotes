eNrtW11vqzgQ/SvIr6WVgXxL+0ATbi9qQlggaaubVUSJ26INkAVy226V/762SSE0uEmbVNrd6z64
YM94PPaZgTkiL0APk9QNPZSAzgsYzzwIOuBlApLn4Daam1Hip34UTvDgBDzjf3IDihPwhK/qTbjC
l7phO1P7ZnA+7OPOCfg2d5OHXncczVP3Hk0AFlnE0QLFqY8SKvHjZTKZgLHaH2nkokOaBmlE0th9
vadZlvb7SLe0Xi5w584TlAsZqqOPtamhDoopRsUUptbV1f50ZOhOWSYX6Wl219JNRx8a+eDPbMmC
Hwpk9cmGtd1myu4UMt+HV1PTGpqa5dzkw2m8LHyxR+dd3eqO2JN813s9zWBsRWkVPe2bOuo7Ff6O
BqZ63td2LqF6uwa68WZxsEpZz84rXM7ndGj7AMZiMBaX41y5Yu9EdAoV0hSYGKjXTPPOjVl0W5ra
L8/9dkeo4uoPistNFBFgYvTTfi8KFlGIwtRwA0RHZt7pGtCndrSMvQzXmyDKpIRXDCWFVByl7jqG
JkCSaJ+/DrrcAAk8OlIRcUrzrP4aczX5rE6iTuvpDj1PokzPsrTwafq8yCZ2Q3ce3dPRZHnbQ4kX
+4t8OSPhN6Eh4OMIqURf72qGrU3pnpJxuO4+t1TrZnphDUcm7c/mQ3PkpWhmlsN7lHmNfQ7vs3jP
dvtu7i/o/Qn+oz25GbrxKyACS943+7QgO/tYKPGTNIr3TT7S4cnHOjT5ZGsmmKhOOxZPOwekneFD
kIiXtB2Q9v38c0Lyz8nX5B+KtZVYgUK5cdaqH45EBwWLQ8GY+MFyTpOWkOLpEA7mZUwfjDN0HyMk
dNHc85eMJyR7BR9C6xu8fRSuZaT9p9D6Hjq/ApNMSMIjwNGTDkXjnR8nqRDFMxSX4OhF6O7O93z8
vGMAkWWb4/AXxKF8cFZEXhTOPgdEmQPx/wDEYz2jwyg4FI2bAHRT4fHB9x6EhRvjiiJFcSI8IjyA
ntLYJe/oDFwy18GB+e8FZnXxajFK11Ix9LZivUAhin1PKAntVbBaMqtcrb+WaM167ajFqoWLVUm4
zN7fj1iwWlsFa9Uj6Aw7xsbf7ph/N5gH7hN+5Q6E2xi5fwqLCAev4HpxlCRCvD6as+oQNrFqGTOl
4eBKvBIvr/aoSVgwpmwMrYneyQJ5iJTwbBI/dpaTq530gLUmB6Qd5ADMkcfJAU4OcHKAkwP8lYOT
A5wc4Djk5AAHIicHODnAyYGjkgMQMsgBiUEOSO3XEq3ByQFODhyTHJAbjcb7/EABvlaNzQ9c+THq
u7doXkkQVIcXI7qKad6GlhHNkFAM7xdUxENWXDWVM+n1I5GWpFSEVraln4it7PiOE00f/zRkvUnk
iC/C2Y6P0xRpn4/TLuJoGc4+cLwXa+ntE96Yait7FkN7HS/xjkWptovvf1qfz5ofO8EPnRLdIRqG
yg6OLmeH2/IROTrISTpO0nGSjpN0vCblJB3HISfpOEnHgchJOg5MTtKxv+BRWOVmLedJml9A0kHO
0v2iLN1KBN1XyCRjHz2CDrC9BxTgc/OACP6OogB0JAhFoP21pAhOQOfHyxs2AWvJbfgkQ6yy8EMn
uoj9Ge6EeB0iIPwd/S1jC0IZwrZMWnKfRteUdRDBXRwF1/QnRCLuvcm+HKK92TVeZ71J1BqNkjK+
zZWxAFMZT6xQy8pOy8qGskKVmzViM1t8rtyChTIWYFrOvCWtVG2ZXmfKUrXPpK0VytTPbZ9rVZbb
7/lcWN70GetkG7b2Wa72eeOo5IplK1RZYWxYsezt3SbetmA2xQ6fS8tuwRXWtvMqu8hHZBb7StPM
qWqo/Rtbt0kPoblUo6tNTdXCwe1oFgYsxm8mqRm9zVssajlbHfSBmvXSqFRxqn3GiQV0SEIWCxMk
e5RnJ3kOW6DxumFzY8ZcmUTs2shQNxybXK9Wq38A8dxItw==