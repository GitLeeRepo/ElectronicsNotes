eNrtXW1zokoW/iuUn5KKk+luaNBU5YMTvVnrRuMS49yp660UgyShViULOC87lf++3c27AqICkglT
UxCBfj1PP6e7Oefwq3GnL1ZzxdaN5cg0XjTT1jWrcfGrcfe51xs9dIadmy93/Tt6pT+8G3eGV72H
8ZdRr3HRaDQbo9v+cHzn/O3fHnXkzqA37snOdSej3rDrJjG+a2Znqcx/WjopyDZXmvcMSS+Pw4nY
hYf7YX+8VsSQFBDNvfPppkdKeFTmlhYq00/8+tpsfNZNp21tBDAE5CjygP5+NI3Fl8YFudZs2MZf
jQtyq8muen/bBrlPnia5YAmIGLQAPYYSk19uYnLLT0we9hJjNzECgB4jJSPgJWYJNhIjr2TMA1Gk
x3C1eS8xuRWTGHuJeUSrTY6hxDxKrza577aZVXutzVuq7bRZwAC2ATlG20yuuYkFHCQWcLTN5DdG
NDEWI21G6YnJ025vS8Bpebi3pfRqO22GEgRCC8AWT0+h5OSXm5ze89PT590MyBM0A3LCALATjFTe
7zbI8vIycDN2kMgyINKSAD0JkX7npSADEM4A+DXAThPagBcBPZFb4QxEPwOpHW5C288A0AxatP2A
HFGkA6HfA61Q/Vt+9RHy2s+3WPuFSPv51rb2C077SffS6m9IIFT9iARafFQCDmDpUYwfqgmwFT35
0+pTGICE6jORx8jf6TxA+WWDZUQ+jmVaYINlyLilRzF+rMdX3cE9JB1EgUNOaz0fAIcPcQV0O9Tv
eaHtjXewfbwLPmhEr92Ez+gRxXNcmGmCdjugoQQFaKfx0T4H6Z3Gh3p8k5r59JJdmmozpmmvtTnE
NO30NqPNgYJQ7EDZbDPGNDGOVBvj9MSYVZv0BxmOGx0WDNF4XeZ0mCRQlNHyEzRKuMPIwxGNQvqA
8nqbcmw8r8d2GHnal/OmOtoCEt7vMKfaeHu11zvMHdCbpCiABFJcG9cuHzNei5Qv4AReW6Nl0pHu
AAHbB0jQ6wh4rOqWjkGm0gOtAlyxOUoxKrZ4pbguNo/THW7MQIpB6XzLoybCMZtKQYDx1d+gJjYV
2CRGMbb6axOCFlPFmyMNpuuzEHCctq/1/FaF4PY8mwJtTv749Kr7kz8CAKKakkATP/lzQONMgeiR
j5/8JUyE+PA8ZqPdoXlMgsxpu0kOV8bixVhqS9ua6Np3Mh2/U5+1BVl0qHRSv7RsZak6M/PuYIDJ
/V/TxuNcf5k2LqaNM/Jv2mhOG6qXy1BZaOxWV3/SbWX+YbCa2/pCszXzA4IAsKdf/NUMe/TXdDpt
3C91m54v6AECbkLPTXpgq5Lgln/9zliZqjb++aL5NyfdK3p6ZaXQFcnD3ZfBp9sbVswfc8V6Jo3w
q2H9XHw15iPD0ukSizxDmvaTnHgyrKeNH1OKcDowpo1hZ9yfOEsbp3GDAcvBNGzFTTttuLl2e3dX
cn807t8Owx3BBR3B+TWIKRtgv2zMyr7pf5I78peHa/n2fsRyjPb4g017gF5XyMrNeGJ3dVdwgTiI
8NgdukCMtOGmf9Ub3jkrR3YDssu9bn9MF27sEl0JOg0mzV0+sWt//0M6mmBkMlNBdljM1A8TY24r
T9oHR35xgPibIWLSubnv+aIVA7nf9Ls9We79+74v97r+A2x56T8Ulpj3xH2Qxah31e/csBVo9Bn/
kbAYvZvfnJpz+pKjjbBCpW0vJtqc4Jl/3X5+GMm3o548/uLfZh3uP3L/6aovX90nZ/KvfrfbGyZ0
RaQW3d4fnfubcUx77wcjJu9tVYjvrkF/uFY5EJe478hruZrP2a1NAUyai0lzFYz+mL5rah8ATw8B
JgadvxKLZ8D2Lsu9zk007/UeYQlf/0mhkCsXwakkgrBHIliK5RAybjY5BMJYDpmpnIc9Kxg1MYUi
6dzjDyygc5wfgdBhHiUQrwEbBOKyqzbXVFubjaJj+z6FXazV165mqab+4nfIPXfJiVQZLJP4R4bZ
2UfWLN2yDTMr6cDDSUc+lHScOlNZxNONXNPNAXRz+7ywmn+y44Ae03nnjPLOWTG8w7D22oxBIRLP
W/hwJI61xcuhYLT8HWnOJtlpZDyuTKYQZ9qTqWnclTZX9VWCZkyuwU5oXcPbrnCNIu1NoTUNnUVg
MhGSIAc4qvBQND7qpmVzhjkjc+owHFVDe3zUVZ1QfwIQk8qucfgOcYgOZkVNNZaz/YCIaiD+DkDM
S0cvjcWhaAwDULG578+6+sy9KKbCNh8s7rtGbmg/bFOh0/MEXCbWowZmdYGZsmiNrHwS16zAW7NK
IHbNKmfe9brWlpqpq1yk3M0S6QsJp0QRC3kuV2UYXazKeyxV5d2WqjJZqkLuT2cVsblcjdNe5wiD
ZOhup4tUHhgoP8hsfcF9NTXlP9wL3UXlFNU0LIszXamcx4/+EUkahVvk9uJz83Pzz88ZljNJI4Bt
4LDlVAqB+KMrMhT83eDUleiruzkwJjwnZN8foI9/6CyXPsCTtgkiVRr3/hond4bfjGgXTC5Fusk1
Xcr8JaSgcX4Ilyj4wZ+R37z/e4IuhUkm8ojDihI0Kw01TuvpAo92Rjw+YrJKIcetpFuI7ogm3zK2
Uml/uxbOpprSMsgyX8iihhPupWkGKuY1yCfpB8nXDxDGb2rGZJZFW3RmM8KTDuLiFYXYDopGOb4X
YQQRVRV+LXbTFrspi6TdzO5gwL+Ll2yCL1BBKvkdm4C9PXJByPcVG1/MKzaKSFRJLUZ010d0Ip6S
0wk8g6fiIbOZgjVUJpKugrLKpA0OVVl7LWbS5hzHV0/Ugs7VEYAvVz1RSxin6HYrZ+2EKqSdaOFS
JYmoqy0M0nukzprFKf7b0pn+TZ9p5jk3fvZenXr3nCk1p1ucODnnuP6Ss5/JD1WxNPKX/xh9QF3Z
9BUH+shztsEJ7JblTslJUpI5eYj8p0Y2LO2jYdL3JJyMPp7IkDsjf5w2aRasCO2HsniZaxcsB0SJ
E51yhknzPw8yW1BdRh6bcd91+zlSpQmtxpP+zamoWxH/rvHoVfG8ZuOajY/FxlgMZuxCuWyMcaAI
2jnTsVQhOp4gJTsZ3yhftXksBafIm7rlBAmTRB3s4rXiJZ1ZtkNjpnFBgTFFSfw59KbvLcjnauKC
lKhwg4ocKl2HLWLF64z0ePF+rYR4qZl9SeLFoEjxfq2UeK+Xsx0WddemsVrOdhVwKNV26UIh3tr1
2s0h075/UGCcdH3jVgG38pQt7cuocL1KJ4h2F/NWWJu31uattXlrdCi3jmDeinGR5q2wmuatOE/z
1n1sEpsF28XmaPSa90IyT55KZ6AyF5CJNq8FLCijNrOu6cwetg3Ncsxiy7R5rdiuRwSO1QFr4bsd
eUIyZ7PYcmxeaxzWOEw3iy3J5rUG4m8HxCLMYsu3ea2BWfX3EpnMW4XAr1uCWe1bE5asGe1bBd4v
UhTzNXDFlTRw3c+Mc6fF529iNZu6WNxqM+sZuMpCBbcH0N5GqrntCuRujvp2tgL2NEZN3BUo0ji1
tO2BXYFY6q5A1WynS5xgVN5yuphl2c5wLGVXoMZhjUNQhV2BGojvA4gH6ujydwVqYL5JH6dM2wM4
sGID5ewOBC/RpZy9X4WjbA6genOgUpsD3cEAvgtnMugb/LZByc5kMDBXlPJ1JoPFOJORfIT3EcYz
2HttwZJRgdq+paPUyhcWQnE+hhC8Bd8eS6feM5yqm+pKtx3vGGM5/8lBl4SJaPZ39zmZoFOSz0Ih
fc+tluqzsnxiPjjPpGhn99vxuPHKOk9x/8EnkyS/H/EEnubk7SOue/vUoQHq0AAle/vQEOEO4SGA
y/X2EUBQNMjZ2weCCrn7XC9nsAIOA6K0xfQ3N38BEQfWvnm7C8Bi3AUoQMRKalHhEn3kqau+63Eq
1uqisu6ghyqNLTqtApFkYOChWbJzaBDEpp23b6hYLWUBKqAsgm8pFK0seFScsgDFKAu6in0fwX5a
R9ufEYSi9mdQcQtxXM2QdYi75GTh44nM05AWwmkdjK6eQhxtCiFKR5tCiGJhUwhcsWg/sAAmimOV
UKCcyeH24tsCzmR/45NHeJsyQybn4hudWIc3FTR5u47LK+4Yf7y4Y6iwuGOwQkwko0o7QacbXtTe
z1WMovVbOkHvDsTa+zkO6+8u5Fsx1qV7wLH2fq5xWAkc1t7PNRCroqNr7+camLl940cs28o5+BJu
3lbOqHaBrq2c2c5Eq+Lf+MGhb/xMkHO5fnNS2+odJzI3DgzmWiVH5haCovmcNyxb1fqMD3gfnhfi
0T7jA1FRn/EBxb3Z5yuuqGD4Y3Qo/AOekd8orMX4WovVWux4X/sJfV9CLPmtW/B9CQhz1mJ8lb4v
MVNRHfu8jn1exz5PCuqW8MWEIoKfCyAIfg4FnHf0c1TJ6OcTpFbiEyihT8tJuOBvoPA49A0UKKGc
P4KiVuojKDKfp2VHgVHq99Qre5py1BrlMCOOrUYYeasWGHprVHyY+j3BWJQtR5kGjlGkvSm05mve
mO11ZCwkcw5Tvyca87flqHH4DnGIDmbF/G05aiC+LSAWEaZ+TzQWa8tRA7O6wDw4fp2/LSFltuxI
crTNGL/O9z4Qc7bs4Ctp2fFbGmFsMTzZaobR3N/mJWklGrbsaFfXFfZExrULbO0Ce0RDjuDTve2S
gy7hIIBHO++gS+2q+cDCSnKQeAlPxNNDFFDBFFRhI+KKO6cd04p4F/4Rj8c/uDj+gbBiBPQmwnJ6
LzFn+jd95oTF3DcGJ722sum+NPyIaPRL3olw6RoekaQpMTdDkQQSQm9CGgANnnKGSfPPKQgnXwfh
rOeDR+ZjFMwHYcmBCFAooFvekQiqE4Pztdn4n2EsaCNBs9H774r1nNW4+PtX40Vfjo1rU58RsgaE
uKNCIhdRG/xAgMj69f8yZEcX